LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;
ENTITY RAM_8_BeachWilliam IS
	PORT(LOAD, CLOCK: IN STD_LOGIC;
		 ADDRESS	: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 D			: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 Q			: OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
END RAM_8_BeachWilliam;

ARCHITECTURE Behavior OF RAM_8_BeachWilliam IS
TYPE RAM_ARRAY IS ARRAY (7 DOWNTO 0) OF STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL RAM_SELECTION: RAM_ARRAY;
BEGIN
	PROCESS(CLOCK)
	BEGIN
		IF RISING_EDGE(CLOCK) THEN
			IF LOAD = '1' THEN
				RAM_SELECTION(to_integer(unsigned(ADDRESS))) <= D;
			END IF;
		END IF;
	END PROCESS;
	Q <= RAM_SELECTION(to_integer(unsigned(ADDRESS)));
END Behavior;